module FD_pipe(
    input wire [15:0] instr, 
    input wire [15:0] next_pc, 
    input wire [15:0] pc_inc,
    output wire [15:0] FD_instr, 
    output wire [15:0] FD_next_pc, 
    output wire [15:0] FD_pc_inc,
); 

//not entirely sure how to do write_data... coming from writeback


endmodule