module MW_pipe(); 

endmodule