/*
   CS/ECE 552 Spring '22
  
   Filename        : fetch.v
   Description     : This is the module for the overall fetch stage of the processor.
*/
`default_nettype none
module fetch ( input clk, 
               input rst, 
               input [15:0]   pc, 
               output [15:0]  next_pc, 
               output [15:0]  instr, 
               output err);

   // TODO: Your code here
   
endmodule
`default_nettype wire
