module DX_pipe(); 

endmodule