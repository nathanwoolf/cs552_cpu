module XM_pipe(); 

endmodule